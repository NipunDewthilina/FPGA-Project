module whole_alu (
    input clk,
    input [16:0] in1,
    input [16:0] in2,
    output [16:0] alu_out
);
ac #(.N(17)) ac (.clk(clk),)     


endmodule)