module instr_mem #(parameter width_in,parameter width_out)(input clk,
// input read_en,
input [width_in-1:0] addr1,
input [width_in-1:0] addr2,// not used
input [width_in-1:0] addr3,// not used
input [width_in-1:0] addr4,// not used
output reg[width_out-1:0] instr_out
);

    reg [width_out-1:0] ram [2047:0];

    localparam ldac = 5'd3;
    localparam nop = 5'd28;
    localparam mvacar = 5'd10;
    localparam mvac = 5'd9;
    localparam mvacr1 = 5'd11;
    localparam mvacr2 = 5'd12;
    localparam mvacr3 = 5'd13;
    localparam mvacr4 = 5'd14;
    localparam mvr1ac = 5'd15;
    localparam mvr2ac = 5'd16;
    localparam mvr3ac = 5'd17;
    localparam mvr4ac = 5'd18;
    localparam ldiac = 5'd5;
    localparam stac = 5'd8;
    localparam add = 5'd19;
    localparam mult = 5'd20;
    localparam lshift = 5'd21;
    localparam sub = 5'd22;
    localparam inac = 5'd23;
    localparam jpnz = 5'd24;
    localparam jmpz = 5'd26;
    localparam endop = 5'd31;
    localparam clac = 5'd30;
    localparam stiac = 5'd26;

    localparam operand = 12'd0;

    localparam nop_addr = {nop,operand};
    localparam add_addr = {add,operand};
    localparam mult_addr = {mult,operand};
    localparam lshift_addr = {lshift,operand};
    localparam mvacar_addr= {mvacar,operand};
    localparam mvac_addr = {mvac,operand};
    localparam mvacr1_addr={mvacr1,operand};
    localparam mvacr2_addr={mvacr2,operand};
    localparam mvacr3_addr={mvacr3,operand};
    localparam mvacr4_addr={mvacr4,operand};
    localparam mvr1ac_addr={mvr1ac,operand};
    localparam mvr2ac_addr={mvr2ac,operand};
    localparam mvr3ac_addr={mvr3ac,operand};
    localparam mvr4ac_addr={mvr4ac,operand};
    localparam sub_addr = {sub,operand};
    localparam endop_addr = {endop,operand};
    localparam inac_addr = {inac,operand};
    localparam ldac_addr = {ldac,operand};
    localparam stac_addr = {stac,operand};
    localparam clac_addr = {clac,operand};

    localparam addr_i = 12'd4094;
    localparam addr_j = 12'd4093;
    localparam addr_k = 12'd4092;

    localparam addr_n = 12'd4091;
    localparam addr_2n = 12'd4090;
    localparam addr_3n = 12'd4089;

    localparam addr_l1 = 12'd2;
    localparam addr_l2 = 12'd72;
    localparam addr_l3 = 12'd91;

    localparam stac_i = {stiac, addr_i};
    localparam stac_j = {stiac, addr_j};
    localparam stac_k = {stiac, addr_k};

    localparam ldiac_i = {ldiac, addr_i};
    localparam ldiac_j = {ldiac, addr_j};
    localparam ldiac_k = {ldiac, addr_k};
    localparam ldiac_n = {ldiac, addr_n};
    localparam ldiac_2n = {ldiac, addr_2n};
    localparam ldiac_3n = {ldiac, addr_3n};

    localparam jpnz_l1 = {jpnz, addr_l1};
    localparam jpnz_l2 = {jpnz, addr_l2};
    localparam jpnz_l3 = {jpnz, addr_l3};

    initial begin
        ram[0 ] = clac_addr;
        ram[1 ] = mvacr1_addr;
        ram[2 ] = ldiac_i; //loop1
        ram[3 ]  = nop_addr;
        ram[4 ]  = nop_addr;
        ram[5 ] = lshift_addr;
        ram[6 ] = nop_addr;
        ram[7 ] = nop_addr;
        ram[8  ] = nop_addr;
        ram[9  ] = mvac_addr;
        ram[10 ] = ldiac_k;
        ram[11 ] = mvacr3_addr;
        ram[ 12]  = nop_addr;
        ram[ 13]  = nop_addr;
        ram[ 14] = add_addr;
        ram[ 15] = mvacar_addr;
        ram[ 16] = ldac_addr;
        ram[ 17]  = nop_addr;
        ram[ 18]  = nop_addr;
        ram[ 19] = mvacr2_addr;
        ram[ 20] = mvr3ac_addr;
        ram[ 21]  = nop_addr;
        ram[ 22]  = nop_addr;
        ram[ 23] = lshift_addr;//21
        ram[ 24] = mvac_addr;//9
        ram[ 25] = ldiac_j;//5
        ram[ 26]  = nop_addr;
        ram[ 27]  = nop_addr;
        ram[ 28] = add_addr;//
        ram[ 29] = mvacar_addr;
        ram[ 30] = ldac_addr;
        ram[ 31]  = nop_addr;
        ram[ 32]  = nop_addr;
        ram[ 33] = mvac_addr;
        ram[ 34] = mvr2ac_addr;
        ram[ 35] = mult_addr;
        ram[ 36] = mvac_addr;
        ram[ 37] = mvr1ac_addr;
        ram[ 38] = add_addr;
        ram[ 39] = mvacr1_addr;
        ram[ 40] = ldiac_k;
        ram[ 41]  = nop_addr;
        ram[ 42]  = nop_addr;
        ram[ 43] = inac_addr;
        ram[ 44] = mvac_addr;
        ram[ 45] = mvacr4_addr;
        ram[ 46] = stac_k;
        ram[ 47]  = nop_addr;
        ram[ 48]  = nop_addr;
        ram[ 49] = ldiac_3n;
        ram[ 50] = sub_addr;
        ram[ 51] = jpnz_l1;
        ram[ 52] = ldiac_i;
        ram[ 53]  = nop_addr;
        ram[ 54]  = nop_addr;
        ram[ 55] = lshift_addr;
        ram[ 56] = mvac_addr;
        ram[ 57] = ldiac_j; 
        ram[ 58]  = nop_addr;
        ram[ 59]  = nop_addr;
        ram[ 60] = add_addr;
        ram[ 61] = mvacar_addr;
        ram[ 62] = mvr1ac_addr;
        ram[ 63] = stac_addr;
        ram[ 64] = clac_addr;
        ram[ 65] = mvacr1_addr;
        ram[ 66]  = nop_addr;
        ram[ 67]  = nop_addr;
        ram[ 68] = ldiac_2n;
        ram[ 69] = stac_k;
        ram[ 70]  = nop_addr;
        ram[ 71]  = nop_addr;
        ram[ 72] = ldiac_j; //loop2
        ram[ 73]  = nop_addr;
        ram[ 74]  = nop_addr;
        ram[ 75] = inac_addr;
        ram[ 76] = stac_j;
        ram[ 77]  = nop_addr;
        ram[ 78]  = nop_addr;
        ram[ 79] = mvac_addr;
        ram[ 80] = ldiac_2n;
        ram[ 81]  = nop_addr;
        ram[ 82]  = nop_addr;
        ram[ 83] = sub_addr;
        ram[ 84] = jpnz_l1;
        ram[ 85] = ldiac_n;
        ram[ 86]  = nop_addr;
        ram[ 87]  = nop_addr;
        ram[ 88] = stac_j;
        ram[ 89]  = nop_addr;
        ram[ 90]  = nop_addr;
        ram[ 91] = ldiac_i; //loop3
        ram[ 92]  = nop_addr;
        ram[ 93]  = nop_addr;
        ram[ 94] = inac_addr;
        ram[ 95] = stac_i;
        ram[ 96]  = nop_addr;
        ram[ 97]  = nop_addr;
        ram[ 98] = mvac_addr;
        ram[ 99] = ldiac_n;
        ram[100]  = nop_addr;
        ram[101]  = nop_addr;
        ram[102] = sub_addr;
        ram[103] = jpnz_l1;
        ram[104] = nop_addr;
        ram[105] = nop_addr;
        ram[106] = nop_addr;
        ram[107] = nop_addr;
        ram[108] = endop_addr;
    end

    always @(posedge clk) begin
        // if (read_en == 1)
            instr_out <= ram[addr1];

    end

endmodule


