module processor #(
    parameters
) (
    port_list
);
    
endmodule